library ieee;
use ieee.std_logic_1164.all;

entity top_level_test is
generic(n: integer:=16);
port(reset,clk,l_p,new_data: in std_logic;
     --input_test : in std_logic_vector(2048*n-1 downto 0);
	  cls_signal : out std_logic_vector(9 downto 0));
end entity;

architecture behav of top_level_test is

component extern_memory is
generic(k: integer:=8;
        n: integer:=16);
port(reset,clk: in std_logic;
     cls_out: out std_logic_vector(9 downto 0);
     q: out std_logic_vector(2048*n-1 downto 0));
end component;

component top_level is
generic(k: integer:=8;
	n: integer:=16);
port(l_p,clk,reset: in std_logic;--l_p=0 => learning process. 
     input_vector: in std_logic_vector(2048*n-1 downto 0);
     input_cls: in std_logic_vector(9 downto 0);
     new_data: in std_logic;
     class: out std_logic_vector(9 downto 0));
end component;


signal q_s,q_s_top: std_logic_vector(2048*n-1 downto 0);
signal cls_out: std_logic_vector(9 downto 0);

begin
u0: extern_memory port map(reset,clk,cls_out,q_s);
u1: top_level port map(l_p,clk,reset,q_s_top,cls_out,new_data,cls_signal);
q_s_top<=q_s when l_p='0' else
         "00000000000001000000000101010010000000011001110000000011101000100000000110011110000000000010110000000101101111000000000100111110000000100001101000000001101101100000000110111110000001100100000000000101010001100000000010110100000000010100111000000000110110000000000011100100000000100100000000000000011101100000000101001110000000100001011000000000011100000000000011100000000000100101011000000100000001100000000001010100000000000100010000001000111110000000000111101000000010000000100000000011101010000000000010011000000000001000000000000000100111000000000010001010000000011001100000000001111001000000000001100100000010000001010000000100010101100000011110111110000000110000110000000011100011100000000000001110000000000000111000000101001010100000000101110000000000011000000000000000000110000000000110110100000000011111100000000000100101000000000000101110000000000001101000000001100110000000000000101100000000000110001000000000101000000000010100111110000000000011100000000001010000000000100111011110000000000001100000000100101111100000001000100010000000100000001000000011011001100000001001011000000000000011000000000011101001000000000101100110000000101001101000000000010010000000011100101100000000101010010000000000001010000000000100010110000000110000111000000010010010100000001010110110000000100001110000000000000100000000001010110000000001110001011000000000011101100000000011001010000000010110011000000000010100100000011100001110000000000000000000000010101111100000000011100100000000010001001000000001001011100000001100100110000000100100111000000001101101000000000011010110000000011110101000000000000000000000000011011000000000011111111000000000100100100000001010110010000000001111100000000000101001100000001101110100000000000010100000000001111001100000010011001010000000101110011000000000111000100000000001011110000000100110000000000010010011000000101010011000000011010000010000000100101011000000011100001100000000000010100000000011111011000000000010000010000001010010001000000101111111100000001101100010000000010011110000000001110001000000010111001110000000011000000000000000010101000000000111010010000000010101101000000011001001100000001000011100000000010101001000000010111001100000000001110000000000101011000000000000011010100000010101010000000000101010100000000011110010100000010000000110000000100000100000000111110011100000000000100100000000011110101000000100110111000000000011010010000000000010110000000000001100100000000000110010000000110111111000000001011110100000000011011000000000110101011000000100011111000000000001110000000001000001011000000001010001000000000000100110000001001100011000000001101101100000001110000000000000110110100000000000001011100000000110001110000000000000111000000100110100100000000000000000000000011001000000000000011110100000000001100010000000000000100000000011010001100000000001010110000001001010000000000000000000000001101001000000000000000010000000000001100000000000001010000110000001001011111000000000001111000000001000110110000001011011011000000001010111100000000001100000000000001101110000000101011010100000000001010010000000010100101000000010011110100000100100100010000000011010100000000010100110100000001000100110000000100010101000000000001101000000000010101010000000111110101000000001000110000000000011101010000000000010110000000000010111100000000111100010000000000110100000000000011011100000000000111010000000010011010000000000000100000000001010011010000000010100010000000010011101000000000010101110000001101010110000000000000001100000010001101010000000001100001000000000110110100000011101000100000000000101010000000010011100000000000011011000000001110000110000000000011101000000000010101010000000011101101000000001010000000000010001010110000000000111001000000000101011000000000001100010000000000010000000000001001110000000000101101100000000011011001000000100100101100000000011101110000000011100000000000000010101000000001011111110000000100000101000000001100011100000100100001010000000001001111000000010000101100000000100110010000000000011000000000001000010000000000001000100000000000110000000000000101101000000000010000110000000000011100000000001010111000000000111111100000000101011101000000011000101100000000101010110000001000010001000000000010111000000000011001010000001000001111000000001011110100000001011101100000000010010000000000001110100000000011000101110000000011101100000000000000010100000000101001110000000001011101000000001011000100000000111011110000000000010011000000010111010100000000110001010000000100100100000000000011110100000000001100000000001110010000000000000001001000000001000000010000001000010111000000000000010100000001011111110000000100110110000000110111100100000010000100100000000100100110000000001000011000000000000110000000010011001111000000000111101000000000011010110000001001000000000000110101000100000000010010100000000011001001000000001011100000000001111101000000000010000000000000000010001000000001000001010000000110111111000000000001000100000000000100100000010001101000000000000100100100000011000111000000000010000001000000010000011000000000111110010000010101101000000000000101001100000000101100000000000100110111000000011010000000000010111010000000000000100010000000000011001100000010100101010000000000110001000000011101101100000000111001010000000110110011000000010100001100000001000011110000000000111111000000001111101000000000001010100000000101111011000000000000000000000001011011110000000010010000000000001011100100000000010001010000000000100010000000000011011100000000010101010000000000000110000000000010111000000001000011010000000000011110000000001001001000000000101101010000000000000000000000000000110100000000000100100000000010000010000000000110000000000000111100110000001000000110000000001001111100000000001011000000000101111000000000000111000100000000111010000000000101001000000000010000111000000000000001110000000000001010000000000001001100000000001110010000000000101000000000000100001000000000000000010000000001100011000000001110101000000000101011000000000101011001000000001101001000000000010001010000000000001010000000001111110100000000000000000000000100100001000000000010110000000000010001010000000000011001000000010111011000000000101000000000000001110110000000001010011100000000000110010000000100100011000000010110000100000000000010000000000101101111000000000010000000000000101000110000001010111110000000000001111000000001100100000000000000000010000000000110100000000010111000110000000010001011000000000100011000000000011011010000000110001000000000010110111100000000100011110000000010111011000000000010100100000010001110100000000011010000000000010011000100000000000011010000000101010010000000001101001000000000000111010000000100110101000000000100100100000000010011100000000000001100000000001101111000000000001010000000000000000110000000011101000000000000000000110000000000001101000000000010100100000001010001000000000001100110000000010110011000000001010110110000000000100010000000001000100100000010001101110000000011000101000000011110101000000000001110010000000001100111000000011001111100000000001001110000000000100001000000000001000100000000100010000000000000100000000000000111100100000000100101110000000000001010000000000111111100000000111001000000000010100100000000001001011100000000111111000000000000010010000000010010110100000000101110110000000010100110000000000011100100000001001101000000000001011001000000000000100000000001001100100000000000110000000000100011010000000101011100100000000011000101000000000100110100000000100101010000000000000010000000011000000000000000001000000000000011100100000000001100001000000000111010110000000001111010000001000000101100000000011000110000000010111010000000001011110100000000000000000000000000101101000000011110101100000000100010110000000000100111000000000001010100000000001101000000000010101000000000000111111100000011001011000000000000000111000000000111000100000000111010010000000000000010000001000111000100000000000110000000000010101100000000001010010000000000010010100000000000110111000000000100101000000000001101110000000000111001000000001100101000000000101111110000000000000100000000001011001100000000011011010000000000010101000000001100110000000000000111110000000001000000000000010100010000000000010110000000001110011011000000000101010100000001100100110000001000101100000000010010100000000000000111010000000001001000000000000010101000000000010000000000000001011100000000000101010100000000011000110000000001110000000000000001011000000000000001110000000000110111000000110010000000000001010100000000000001110110000000001010000100000000110010110000001101010011000000000110111100000000101000000000001001000110000000001001111100000000000000010000000110111100000000001101110100000000110011100000000000001111000000000100111100000000011100000000000010000100000000101111010000000000000111000000000000100100000000000101001100000000101000010000000110001100000000011001001000000000000000100000001000001111000000000110011100000000000001000000000000100000000000011100101100000000000000000000000000101101000000001110110000000000100001010000000001101110000000000101111100000000000000000000000000101111000000011010000000000010111010100000000100100101000000000000001100000000011110010000000011010110000000000000100100000001001101010000000000111011000000000001000000000000001101100000000001010000000000001101010100000000000000000000000000000100000000001011101000000000000000010000000011010010000000010100001100000001000000100000000001001010000000000111101100000000110010010000000011000111000000000010010000000000110100000000000001111110000000001111111100000000001000100000000011011100000000010011011100000000110100010000000000111001000000001111010000000000010101010000000000011111000000001010111000000000000011100000000110011000000000000100000000000000010110010000000010100010000000000000111100000001000100100000000010111000000000000110011000000000000110110000000000000001000000000110011000000000010101110000000000110001000000001101100100000001110100010000000110111111000000001100010000000001010011010000000001101010000000000011101100000011111011000000001011110010000000001100101000000001010101110000000001110101000000010011110100000010000101110000001001011101000000111110000100000001000001010000000001000110000000100001100000000000110100100000010000111111000000000110001100000000000010100000000011011101000000000000101000000000100011100000000001000101000000101011000100000000000010100000000101001100000000000111011100000000110001110000001110001100000000010101101100000010000001000000000000101111000000011010100000000000010010000000000000111110000000101111010000000001111000010000000000100001000000000101101100000001100001000000000010101110000001010001000100000000011011010000000010001111000000000011011100000000010101010000000001101001000000000001000100000000001011000000000001001111000000000110011000000000010011110000000000000100000000001010011000000000010000010000000000110011000000000011110100000000010000100000000010001100000000001100101000000000101100110000000011001000000000000011010000000000000100010000000001100101000000001001100000000000000110010000000010000111000000001001110000000000010101110000000010011100000000001101011000000001000001010000000011100100000000001000001100000000000111110000000111110011000000000100100100000000011010100000000000010011000000000010101000000001100011010000000000000000000000010001111000000001000011110000000001000100000000000100001000000000001011010000000011111010000000000110100000000000010011100000000001001111000000001000001000000000000011000000000110001011000001000100101100000000000101000000000000001100000000000111011100000000000000000000000101010001000000001000000100000000111110000000000011010110000000000110001100000000001100000000000011100011000000001111010100000000011100110000000000010001000000000000000000000000001111010000000001001110000000000001000000000000010111110000000000110000000000000101011000000000000000010000000111110001000000010110000000000000100100010000000001101100000000000011010000000000000011110000000000100111000000000000100100000000101000100000000001101100000000001010010000000001001011110000000100101010000000001011111100000001000110010000000000101001000000001011100100000010010000010000000000011101000000001100101100000000001111110000001010000111000000001011000000000000010000100000000110001011000000001101100100000000101111010000000011001101000000010010100100000001010000000000000111000000000000001000010000000010000011100000000000101100000000011001011100000000111100110000000111000011000000010011000000000000000001110000001110010110000000000100110000000000000100110000000000101111000000000100010100000000110000110000000000000000000000000011100100000010111001110000000001111100000000010100011100000000101011100000000001000010000000001000110000000000101110110000000010111101000000000011100100000000000100010000000001011111000000001001000000000000001011000000000001001100000000000010001000000000100101110000000110101000000000001101100000000001001110110000000011011001000000001111001000000000110000100000000101001000000000011101011000000001000100110000000101111000000000001011101000000000100010110000000000100100000000001100011100000001000010110000000001001101000000010000100000000000101011110000000001101010000000000101111100000000110010100000000000010010000000001000110000000000101001010000000010001011000000001001001100000000101011100000000000001111000000000010110100000000011000110000000011011100000000001101001000000000111000100000000001001110000000010110010000000000000001110000000000101010000000000011001100000000000110000000000010000111000000010000010000000000100111010000000001011000000001011111100000000000001101100000000110000010000000010011000100000000111110000000000010011111000000011101000100000000000000100000000111100000000000010110111000000000110100100000000001011110000000000001001000000010000101100000000001101100000000010111100100000000100001010000000010011011000000000001010100000000001101010000000010001100000000001000111000000001001111100000000000110000000000001010111100000011100011100000001000000110000000000000110000000000001111010000000010010011000000001101111100000000100110100000000000010100000000010100010000000000100001100000000001111001000000000010010000000001000111110000000001011111000000111100011000000000010110000000000010010001000000011011110000000000011110010000000010101111000000000000000000000010000010000000000010000110000000000100011100000001000000100000000000111100000000001010000100000000000100100000000000010110000000010110111000000000001110010000000000101110000000001101011000000001110010010000000001100000000000001101011100000001100111010000000011110111000000001000011000000000010001000000000001100110000000000100111100000000000111010000000000101001000000001000010100000010110010010000000010000000000000011101111100000000000001010000001001100010000000100010000000000000100010110000000000100101000000000000100100000001101100110000000011010101000000001110010100000000011110010000000011111001000000010100101000000000110101100000000010001100000000100101010000000001010010010000000000011111000000011111000000000000110110100000000001001100000000010010111000000000010110100000000001000010000000001001100000000000001001100000000000100001000000000110101000000001011111110000000010101001000000000101101000000000000001010000000000110100000000001110001000000111010100010000000000001101000000001000011100000001001100010000000001111011000000000011010100000000110101010000001000101000000000010010000000000000101001100000001000010101000000011100100100000000000000000000000000001011000000000111000000000000001100000000000000001101000000010011010000000000100000010000000000001011000000000011111000000001000110010000000000000101000000000001011100000011101010000000000010011111000000000001010000000001010110110000000000010010000000011001010000000000100001010000000101111110000000011100110000000000110110110000000001110000000000000101111000000001001111100000000001111000000000000010010100000000100011010000000110101111000000000100110100000000000111010000000001110011000000000101101100000000001100110000000001001010000000001100101000000000111111000000000110111011000000001001100100000010000011010000000010010101000000001010010100000000000011000000000000101101000000000010100000000000101100100000000001001101000000000000001100000000110111000000000111000110000000100100000000000001000100000000000011010111000000000010011100000000100001100000000000001001000000001000011000000001001001000000000000101001000000000001001100000000010110010000000010100111000000000011110100000000000100000000000000001110000000000010100100000000010110010000000010000011000000011001001100000010011010010000000110000010000000000001010100000001110011100000000001011010000000000101010000000000001011110000000000000000000000000011011100000000000000100000000000100100000000101001010000000000101010010000000011001110000000000101001000000000011000110000000000001110000000001000011100000011000101010000000001010011000000000001100000000000001010110000000001101000000000010000001000000010001101010000000000101011000000000100010100000001000110100000000001001000000000011010111100000000100001110000000010000101000000000100000100000000010000010000000000001110000000110100110100000000010111100000000000010100000000000000000000000000100101000000000100111111000000001001111000000000001111110000000000000100000000000010111000000000001001100000000011001111000000010011011100000000101110010000000001001100000000000011011100000000010100000000000011000111000000001100101100000000011110110000000001111110000000000010010100000000010111010000000010000110000000000010010100000010111101100000000000101001000000001000010100000010010100100000001010000000000000100000111000000000000010100000000000001010000000000011101100000000000110010000000000110110000000001001001100000000011101000000001011001110000000011101000100000010110011010000000001101001000000010100101000000110000000000000000000100100000000000011000100000010101111010000001010111110000000100010101000000000101000000000000000010111000000101000100100000000000000000000000110011001000000000000011000000000000000110000000001010011000010111010100000000010001111010000000101010000000000111101010000000000011101000000000000001000000000000011100100000000001000000000000101010100000000000010000100000011001101100000000000010001000001001000001100000000010010010000001000010110000000000110011000000000000010110000000000000000000000010010111000000000000001000000000011101101000000000110010100000000000000000000000100010111000000000110110100000000100011100000000110001011000000100110100100000010110011010000000000001010000000000011010000000000000000000000011001111100000000000000000000000000001000010000000000000111000000001110001100000000100011100000000000101000000000010101010000000000000010000000000100001011000000000101011000000000000110010000001000001110000000011110011100000001000000100000000010110010000000010011011100000001101100100000001100101001000000100101111100000001101000010000000110000011000000000100010000000001110001110000000011011101000000101110011100000010101000010000000000010001000000010100001100000000110110000000000000010101000000101110000100000000000010100000000001000001000000001101101100000010010101100000000100001001000000101010101100000000001100110000000011111001000000000000000100000000000000010000001001000011000000001000010000000001010000010000000011010100000000001010101000000001110010000000000010010010000000000011010100000010110101100000010110011110000000011000101000000001000001000000000001010011000000001001111100000001000010010000000000000011000000000110101100000000001010100000001000000100000000100100101000000001010101110000001010100000000000000000001100000000111111100000000000001011000000000001000100000000001110010000000110000000000000011101100100000000010110000000000010000000000000000000000100000000000000100000010000110101000000000001111000000000100111100000000011011101000000010100100100000000000110100000000001001010000000111110110000000001101010000000000011100110000000110111010000000000000000000000000100111011000000001111011000000000011010010000000000011110000000001010001100000000000001010000000011011011000000100110111000000000000000000000000001010000000000110100001000000000000001010000000011101001000000000110101100000000000111000000000101010000000000001001110100000000011111000000000111001010000000001001011000000001000010010000010110100100000000000000000000000011100001010000000101110111000000011000001100000000110101000000000000001000000000000000111000000000011000110000000100101010000000000010110100000000000001110000000111001100000000001101011000000000000111100000000000000101000000000010011000000000001111010000000100110010000000000000010000000101000111010000000001011101000000010110000100000000001100100000000000011101000000001000111100000000110011100000000000100110000000001111000000000000010000110000000001011101000000100110111100000000001100100000000011011000000000000000000000000000001101000000000000010011000000000111100000000000100111110000000000000010000000000001110100000000011101010000000000111101000000101010010100000000000000000000001010110000000000001101111100000001100000110000000101100100000000101101101000000011100001000000000100010010000000000100101000000000001000000000000001100001000000000111010100000000011011110000000001110010000000011011011100000000010000010000000011011001000000000110111100000101100100010000000110010010000000001000001100000000000110110000000000000011000000000111111100000000000100100000000001110110000000000111001000000000000000110000000010011010000000000111100000000001110011110000001111000110000000001110000100000000000100110000001001001000000000010010100100000001101101000000001011011110000000000001111000000000000000110000000010101001000000100001000000000000011000110000010010101100000000010010010000000000001000110000000111000001000000111011010000000011111001000000000000011111000000001110010100000000100110110000001001011000000000000010000100000010010000110000000111110010000000100110010100000000011101110000011001101110000000001010010100000000000110010000000000001011000000001011010100000010101111100000000000010001000000000000001000000000000001000000000000000001000000010010111000000010110010010000000011010011000000000110011100000001011101010000000100000101000000010100011100000000011010100000000000001100000000010010000100000000001000110000000110100101000000101011010100000011110100110000000011011101000000001010001000000000000000000000000001010011000000000100100100000000001000110000000110000101000000001110000000000011100110100000001000010000000000100010000100000000001101000000000000100011000000001101100000000000001101010000000001010100000000000000110000000000000010100000000000010101000000001001100000000000010010000000010011111010000000000100011000000001011101110000001000011010000000000100110000000011001110010000001100001001000001011000110000000001100101110000000100110000000000000011100000000000001000000000000100111000000000001001101000001101001101110000000010001011000000000010001100000000111110110000000110011000000000000101101100000000001110010000000001101011000000011010000100000000111000010000000110110111000000011000001100000011001001100000000111111000000000000101100000000000000000010000000001011111000000011011101000000001011100010000000011111101000000000000101000000000011111100000001000001011000001011101001000000000000110110000000000011101000000010110000100000000101000000000000010110000000000000110100000000001011011010000000111111000000000001111110100000000100001110000000100101001000000000000110100000000101001110000000011111000000000001000101100000000001100100000000001101100000000100001111000000000010110110000000001101010000000000001111000000010001111010000000010001111000000101010111100000000011111110000000011100100000000000011111000000010001000000000010100101100000001010110110000000000000000000000010110011000000000000000000000000000110010000000001001101110000000001111100000000111001100100000000111000110000000010111000100000001100110110000000000000000000000000011011000000001000100010000000111100000000000001101101100000000011011110000000000101000000000000001001100000000000100110000000000001111000000000000000000000011111111110000000000001011000000000010101000000000000000100000000011001011000000101010111100000000000011010000000011101001000000010000010000000000010001000000000010100010000000000000000000000000010010010000000000010010000000000000100100000000001011010000000000100111000000000011100100000000110011100000001101011110000000000001110000000000001111010000001010010011000000000000000000000000000110100000100010011110000000001000001000000010110001100000000001000111000000010001111100000000001100100000000000001000000000000000100000000001000101100000010110010000000000000001110100000011000111110000000000100001000000000000111100000000110001010000000011100000000000000110110000000100011011100000000000010100000000010010100000000010100111010000000000000000000000010101110000000001100001010000000000001110000000100001011100000000000001000000000010101101000000000010010100000000000000000000000001100011000000000000001000000000111001110000001100000010000000001101010000000011000101110000000010010101000000000000101000000001100100010000000000000000000000000000010100000001101001000000001001011101000000001111111100000000000000110000000000000001000000000000101100000011001110110000001001101011000000000110010000000000001000110000000001111011000000000011010000000001011110110000001101000101000000010010010100000000000010010000000000000111000000001010000100000000001000110000000100000100000000001000010100000000000100100000000000111111000000011001100100000001000001100000000001010000000000000110110000000000010000010000001001110100000000000111000000000000100010010000000010011001000000000000001000000001110100110000010011000100000000100000101000000000110101110000000100110111000000000000011100000000010111010000000011110110000000111101011100000000000000000000000011001111000000000110110100000100010010100000000000000010000000010011001100000011100011100000000100000101000000111011001000000000000010100000000011111100000000000101110000000011010001000000000011110000000000000111001100000000000000100000000011011010000000111011110100000001111011010000001110110000000000000100111100000000000000000000000010110001000001111000100000000010100000010000000000000100000000101011110000000000011100010000001000111001000000010011010000000110001011010000000101110101000000010000100100000000000000000000000100010100000000001011110000000000000110100000001001010100000000010101001000000000000000010000010000001100000000000000000000000001011011110000000000000011000000101000110100000001001010010000000001000001000000000000000100000001000101010000001011010010000000110001011100000000001110010000000010001100000000001101110100000000110101110000000010101010000000000010101000000000000001110000000001001011000001100010111000000001001000100000001111001010000000000000000000000000000001010000000000100010000000011001001100000001111010100000001101010110000000010010101000000000000010110000000000001111000000000000000000000000000010110000001101101000000000001001000100000000000110000000001000110010000000000000000000000000000001000000000000000110000000000010000100000000011100000000000101000100000000001011100100000000010111010000000000111110000000000101110100000000000111100000000010010110000000010101100100000100100001000000000000000110000000000000010000000000111011100000000000100100000000000101111100000000000010010000001001100101000000111111001000000011101011110000000000110101000000010110100100000000110000000000000010000101000000001010111000000000000011100000000101110110000000000101010100000000000010010000000100010010000000000111010100000100100110100000001010101010000000010000000000000001000011010000000000011101000011000011100100000000010110110000000000011011000000000000010000000100100010010000000000000110000000000111000100000010101011000000000101010010000000000100000000000000011011100000000001100101000000000011100000000000000101010000001101010100000000000000000100000000011110110000000010010101000000000000111000000000010110010000000100110000000000101101000100000000010000010000000000011011000000001010100100000000001110110000000000001100000000000010100000000000100000010000000000000011000000000100110100000000010111010000000011101011000001001111010000000000000000000000000000110001000000100001101000000001101000000000000001101000000000000000010100000100011101100000000101100010000000000001110000000000000000000000000001101010000000000010111000000000000100110000000110010010000000100101100000000001110010100000000000011100000000010101100000001100101100000000000001101110000000010100000100000000001111000000000000000011000000000100110000000000101100000000000001001111000000011110101000000000000011110000000101001100000000010010111000000000001000000000000101110101000000001110101100000001011110110000001100111011000000000000000000000000000000000000000000111100000000001101101100000000001001100000001001001011000000111110110100000000000010110000000010001011000000000001001000000011000011000000000011100011000000000000101100000010010110010000001101011111000000000000000100000000000100010000000001110001000000011101100100000000000010100000000110011011000000100111100000000100011100010000000010011010000000100000110000000000111001000000000000000011000000101001010000000000011010000000000000000011000000000111011100000000000111110000000111011000000000001100000100000001001100100000000101001110000000000111101100000010000010010000000000000000000000000010111100000000001110110000000000001111000000000100000100001001001111100000001001000111000000000100001100000000110100110000000010111000000000101000100100000000000000000000000010000010000000001000000100000000000100100000001000000101000000101101001100000000100011000000000010010010000000000000000000000000110000100000001000100110000000010011111100000000110010110000010010011101000000001101111100000000010001010000000100001000000000000000000000000000011111110000000111110011000000100010011000000010000110110000000100000000000000001000100000000000001011000000000010011110000000011000100000000000001011100000000100000000000000001000011000000000101110110000000011000011000000010101000000000000010100010000000000011001000000000001100000000010011010010000000011001111000000000001001100000001111000110000000011001010000000101001011000000010000001000000000110100101000000111010100100000000000110100000000110001101000000001100100100000001010000010000000110100010000000000110101100000001101101110000000100100010000000001011011000000000001011010000000010000010000000001100111000000010101111110000000000010110000000011001101100000000000101010000001101111011000000000011011000000000000000000000001101001001000000001001110000000000000100100000000010001100000001000001000000000000000010000000000101111111000000110111111100000001000011000000000001101111000000111100000000000000101000100000000010100110000000010000101000000000100011010000000111000110000000011100101100000000111001100000001000100001000000101111110100000001110100010000000101010110000000001100111100000001100011000000000100101000000000010001101000000000011010010000000000000100000000001010101000000001000001100000000010000011000000000001101000000001100010000000010000110010000000100010000000000001110101110000000101100101000000011100011100000000011001000000001000101001000000011100111100000000001010010000000000000000000000010100111000000001011100000000000000001101000000000101101100000001010010010000000000100101000000010111101000000000101101010000001001000101000000010011101100000000000100010000000000000001000000000100101000000010010011100000001001111101000000000000001100000001001100110000000001111010000000011111000100000001110011000000000010011111000000000101001000000001000011000000001001010011000000000100011000000011101000110000000001000011000000011011101000000000000000000000001010111010000000011111000000000000001100100000001000000011000000000011011000000011000111010000000110111101000000000100111100000000110110000000000010101000000000111001100000000000010111110000000100001000000000001000000100000001110111100000000000001100000000010000000000000000000011110000000001100011000000000000100100000001101011000000000011101010000000000010011100000001010110000000000110010010000000001101101000000000111100100000000000011111000000001101001100000000001110100000000011010000000000001001001100000010001101100000000001001001000000100001001100000000101111110000000001010100000000000110011000000000001001000000000001101101000000000000000100000000101000010000001010101100000000011000100000000011111101110000000000101110000000001101011100000000101001100000000111111001000000000100010000000001101100100000001100101100000000101110101100000001110000110000000011001010000000010001111000000000111000110000000110011001000000000010110000000000101010110000000001100011000000101011101000000001111000100000000000111110000000111001000000000000101010110000000011010100000000001001000100000010000111000000001000011111000000000101000000000010101110110";
end behav;
